module EX_tb();


